`timescale 1ns/10ps

module controller2A(

    input clk,

    input reset,

    output [5:0] w_out,

    output cnt_out,
    output load_w_out,
    output [5:0] b_out,
    output [5:0] s_out,
    output [4:0] ps_out,
    output [4:0] ns_out

    
);

logic [5:0] w;
assign w_out = w;

logic cnt;
assign cnt_out = cnt;

logic load_w;
assign load_w_out = load_w;

logic [5:0] b;
assign b_out = b;

logic [5:0] s;
assign s_out = s;

logic [4:0] ps;
assign ps_out = ps;

logic [4:0] ns;
assign ns_out = ns;

always_ff @(posedge clk)
begin

    if (reset) b <= #1 6'b0;

    else if (cnt) b <= #1 b + 1;

end

assign s = w + b;

always_ff @(posedge clk)
begin
    if (reset) w <= #1 6'b0;
    else if (load_w) w <= #1 s;
end

always_ff @(posedge clk)
begin 
    if (reset) ps <= 5'b0;
    else ps <= ns;
end

parameter T0 = 0;
parameter T1 = 1;
parameter T2 = 2;
parameter T3 = 3;
parameter T4 = 4;
parameter T5 = 5;
parameter T6 = 6;
parameter T7 = 7;
parameter T8 = 8;
parameter T9 = 9;
parameter T10 = 10;
parameter T11 = 11;


always_comb
begin
    ns = 0;
    cnt = 0;
    load_w = 0;
    case (ps)
        T0:
        begin
            cnt = 1;
            load_w = 1;
            ns = T1;
        end
        T1:
        begin
            cnt = 1;
            load_w = 1;
            ns = T2;
        end
        T2:
        begin
            cnt = 1;
            load_w = 1;
            ns = T3;
        end
        T3:
        begin
            cnt = 1;
            load_w = 1;
            ns = T4;
        end
        T4:
        begin
            cnt = 1;
            load_w = 1;
            ns = T5;
        end
        T5:
        begin
            cnt = 1;
            load_w = 1;
            ns = T6;
        end
        T6:
        begin
            cnt = 1;
            load_w = 1;
            ns = T7;
        end
        T7:
        begin
            cnt = 1;
            load_w = 1;
            ns = T8;
        end
        T8:
        begin
            cnt = 1;
            load_w = 1;
            ns = T9;
        end
        T9:
        begin
            cnt = 1;
            load_w = 1;
            ns = T10;
        end
        T10:
        begin
            load_w = 1;
            ns = T11;
        end
        T11:
        begin
            ns = T11;
        end
    endcase
end

endmodule
        